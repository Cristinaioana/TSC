library verilog;
use verilog.vl_types.all;
entity instr_register_pkg_sv_unit is
end instr_register_pkg_sv_unit;
